library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity transmitter_435 is
    port (
    );
end entity;

architecture rtl of transmitter_435 is
begin
end architecture;
