library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity altimeter is
    port (
    );
end entity;

architecture rtl of altimeter is
begin
end architecture;
