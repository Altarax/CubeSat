library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity temp_hum_sensor_int is
    port (
    );
end entity;

architecture rtl of temp_hum_sensor_int is
begin
end architecture;
