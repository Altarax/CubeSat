library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity one_wire is
    port (
    );
end entity;

architecture rtl of one_wire is
begin
end architecture;
