library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity distance_sensor is
    port (
    );
end entity;

architecture rtl of distance_sensor is
begin
end architecture;
