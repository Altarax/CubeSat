library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity top_level is
    port (
        clk : in std_logic
    );
end entity;

architecture rtl of top_level is
begin
end architecture;
