library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity temp_hum_sensor_ex is
    port (
    );
end entity;

architecture rtl of temp_hum_sensor_ex is
begin
end architecture;
