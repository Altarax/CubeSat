library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity spi is
    port (
    );
end entity;

architecture rtl of spi is
begin
end architecture;
