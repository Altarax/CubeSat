library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity i2c is
    port (
    );
end entity;

architecture rtl of i2c is
begin
end architecture;
