library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity uv_sensor is
    port (
    );
end entity;

architecture rtl of uv_sensor is
begin
end architecture;
